module engine

pub fn test() {
	println('hi')
}