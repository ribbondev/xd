module main

import engine
import raylib

fn main() {
	engine.test()
	raylib.init_window(640, 480, "hello world")
}
